/** 
    Aquí generaremos el testbench general para tods y cada uno de los módulos 
**/
module testbench();

    

endmodule
