module tb_shift_register();
    
endmodule
