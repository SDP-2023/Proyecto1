module testbench();

    

endmodule
